module Control( opcode, funct, RegDst, Jump, Branch, MemRead, MemtoReg, ALUOp, MemWrite, ALUSrc, RegWrite);

	input [5:0] opcode;
	input [6:0] funct;

	//Use reg for behavioral
	output reg [1:0] RegDst;
	output reg [1:0] Jump;
	output reg Branch;
	output reg MemRead;
	output reg [1:0] MemtoReg;
	output reg [2:0] ALUOp;
	output reg MemWrite;
	output reg ALUSrc;
	output reg RegWrite;

	always @(*) 
	begin //R formmat 000000  is default
		RegDst		<= 2'b01;
		Jump		<= 2'b00;
		Branch		<= 1'b0;
		MemRead		<= 1'b0;
		MemtoReg	<= 2'b00;
		ALUOp		<= 3'b001; 
		MemWrite	<= 1'b0;
		ALUSrc		<= 1'b0;	
		RegWrite	<= 1'b1;

		casex (opcode)
			/* R format */
			6'b000000: //R 
			begin	
				if (funct = 6'b001000) Jump <= 2'b10; //jr
			end
			
			/* J format */
			6'b000010: // j
			begin	
				//RegDst		<= 2'b10;
				Jump		<= 2'b01; //@
				//Branch		<= 1'b0;
				MemRead		<= 1'b0;
				//MemtoReg	<= 2'b10;
				ALUOp		<= 3'b111; //@ 
				MemWrite	<= 1'b0; //@
				//ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b0;
			end
			
			6'b00001x: // jal
			begin	
				RegDst		<= 2'b10; //@
				Jump		<= 2'b01; //@
				//Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; //@
				ALUOp		<= 3'b111; //@ 
				MemWrite	<= 1'b0; 
				//ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
			/* I format */
			6'b001000: // addi
			begin	
				RegDst		<= 2'b10; 
				Jump		<= 2'b01; 
				Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; 
				ALUOp		<= 3'b000; //@
				MemWrite	<= 1'b0; 
				ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
			6'b001100: // andi
			begin	
				RegDst		<= 2'b10; 
				Jump		<= 2'b01; 
				Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; 
				ALUOp		<= 3'b010; //@ 
				MemWrite	<= 1'b0; 
				ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
			6'b001101: // ori
			begin	
				RegDst		<= 2'b10; 
				Jump		<= 2'b01; 
				Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; 
				ALUOp		<= 3'b011; /@ 
				MemWrite	<= 1'b0; 
				ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
			6'b000100: // beq
			begin	
				RegDst		<= 2'b10; 
				Jump		<= 2'b01; 
				Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; 
				ALUOp		<= 3'b100; //@ 
				MemWrite	<= 1'b0; 
				ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
			6'b000101: // bne
			begin	
				RegDst		<= 2'b10; 
				Jump		<= 2'b01; 
				Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; 
				ALUOp		<= 3'b101; //@
				MemWrite	<= 1'b0; 
				ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
			6'b100011: // lw
			begin	
				RegDst		<= 2'b10; 
				Jump		<= 2'b01; 
				Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; 
				ALUOp		<= 3'b000; //@ 
				MemWrite	<= 1'b0; 
				ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
			6'b101011: // sw
			begin	
				RegDst		<= 2'b10; 
				Jump		<= 2'b01; 
				Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; 
				ALUOp		<= 3'b000; //@ 
				MemWrite	<= 1'b0; 
				ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
			6'b001010: // slti
			begin	
				RegDst		<= 2'b10; 
				Jump		<= 2'b01; 
				Branch		<= 1'b0;
				MemRead		<= 1'b0;
				MemtoReg	<= 2'b10; 
				ALUOp		<= 3'b110; //@ 
				MemWrite	<= 1'b0; 
				ALUSrc		<= 1'b0;	
				RegWrite	<= 1'b1;
			end
			
		endcase
	end

endmodule
