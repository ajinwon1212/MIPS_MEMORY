module Data_memory(CLK, RESET, Address, Write_Data, MemWrite, MemRead, Read_data); 

	input CLK, RESET;
	input [31:0] Address; 	// Input Address 
	input signed [31:0] Write_Data; // Data that needs to be written into the address 
	input MemWrite; 		// Control signal for memory write 
	input MemRead; 			// Control signal for memory read 

	output reg signed [31:0] Read_data; // Contents of memory location at Address

      	reg 	[31:0] 	Data_memory[0:127];

	assign Read_data = (MemRead == 1'b1) ? Data_memory[Address>>2] : 31'd0;

   	always 	@(posedge RESET or posedge CLK) // When a signal is received from control, the process starts.
		if (RESET)
		begin
			Data_memory[0]  <= 32'd0; 
			Data_memory[1]  <= 32'd0; 
			Data_memory[2]  <= 32'd0; 
			Data_memory[3]  <= 32'd0; 
			Data_memory[4]  <= 32'd0; 
			Data_memory[5]  <= 32'd0; 
			Data_memory[6]  <= 32'd0; 
			Data_memory[7]  <= 32'd0; 
			Data_memory[8]  <= 32'd0; 
			Data_memory[9]  <= 32'd0; 
			Data_memory[10] <= 32'd0; 
			Data_memory[11] <= 32'd0; 
			Data_memory[12] <= 32'd0; 
			Data_memory[13] <= 32'd0; 
			Data_memory[14] <= 32'd0; 
			Data_memory[15] <= 32'd0; 
			Data_memory[16] <= 32'd0; 
			Data_memory[17] <= 32'd0; 
			Data_memory[18] <= 32'd0; 
			Data_memory[19] <= 32'd0; 
			Data_memory[20] <= 32'd0; 
			Data_memory[21] <= 32'd0; 
			Data_memory[22] <= 32'd0; 
			Data_memory[23] <= 32'd0; 
			Data_memory[24] <= 32'd0; 
			Data_memory[25] <= 32'd0; 
			Data_memory[26] <= 32'd0; 
			Data_memory[27] <= 32'd0; 
			Data_memory[28] <= 32'd0; 
			Data_memory[29] <= 32'd0; 
			Data_memory[30] <= 32'd0; 
			Data_memory[31] <= 32'd0; 
			Data_memory[32] <= 32'd0; 
			Data_memory[33] <= 32'd0; 
			Data_memory[34] <= 32'd0; 
			Data_memory[35] <= 32'd0; 
			Data_memory[36] <= 32'd0; 
			Data_memory[37] <= 32'd0; 
			Data_memory[38] <= 32'd0; 
			Data_memory[39] <= 32'd0; 
			Data_memory[40] <= 32'd0; 
			Data_memory[41] <= 32'd0; 
			Data_memory[42] <= 32'd0; 
			Data_memory[43] <= 32'd0; 
			Data_memory[44] <= 32'd0; 
			Data_memory[45] <= 32'd0; 
			Data_memory[46] <= 32'd0; 
			Data_memory[47] <= 32'd0; 
			Data_memory[48] <= 32'd0; 
			Data_memory[49] <= 32'd0; 
			Data_memory[50] <= 32'd0; 
			Data_memory[51] <= 32'd0; 
			Data_memory[52] <= 32'd0; 
			Data_memory[53] <= 32'd0; 
			Data_memory[54] <= 32'd0; 
			Data_memory[55] <= 32'd0; 
			Data_memory[56] <= 32'd0; 
			Data_memory[57] <= 32'd0; 
			Data_memory[58] <= 32'd0; 
			Data_memory[59] <= 32'd0; 
			Data_memory[60] <= 32'd0; 
			Data_memory[61] <= 32'd0; 
			Data_memory[62] <= 32'd0; 
			Data_memory[63] <= 32'd0; 
			Data_memory[64] <= 32'd0; 
			Data_memory[65] <= 32'd0; 
			Data_memory[66] <= 32'd0; 
			Data_memory[67] <= 32'd0; 
			Data_memory[68] <= 32'd0; 
			Data_memory[69] <= 32'd0; 
			Data_memory[70] <= 32'd0; 
			Data_memory[71] <= 32'd0; 
			Data_memory[72] <= 32'd0; 
			Data_memory[73] <= 32'd0; 
			Data_memory[74] <= 32'd0; 
			Data_memory[75] <= 32'd0; 
			Data_memory[76] <= 32'd0; 
			Data_memory[77] <= 32'd0; 
			Data_memory[78] <= 32'd0; 
			Data_memory[79] <= 32'd0; 
			Data_memory[80] <= 32'd0; 
			Data_memory[81] <= 32'd0; 
			Data_memory[82] <= 32'd0; 
			Data_memory[83] <= 32'd0; 
			Data_memory[84] <= 32'd0; 
			Data_memory[85] <= 32'd0; 
			Data_memory[86] <= 32'd0; 
			Data_memory[87] <= 32'd0; 
			Data_memory[88] <= 32'd0; 
			Data_memory[89] <= 32'd0; 
			Data_memory[90] <= 32'd0; 
			Data_memory[91] <= 32'd0; 
			Data_memory[92] <= 32'd0; 
			Data_memory[93] <= 32'd0; 
			Data_memory[94] <= 32'd0; 
			Data_memory[95] <= 32'd0; 
			Data_memory[96] <= 32'd0; 
			Data_memory[97] <= 32'd0; 
			Data_memory[98] <= 32'd0; 
			Data_memory[99] <= 32'd0; 
			Data_memory[100] <= 32'd0; 
			Data_memory[101] <= 32'd0; 
			Data_memory[102] <= 32'd0; 
			Data_memory[103] <= 32'd0; 
			Data_memory[104] <= 32'd0; 
			Data_memory[105] <= 32'd0; 
			Data_memory[106] <= 32'd0; 
			Data_memory[107] <= 32'd0; 
			Data_memory[108] <= 32'd0; 
			Data_memory[109] <= 32'd0; 
			Data_memory[110] <= 32'd0; 
			Data_memory[111] <= 32'd0; 
			Data_memory[112] <= 32'd0; 
			Data_memory[113] <= 32'd0; 
			Data_memory[114] <= 32'd0; 
			Data_memory[115] <= 32'd0; 
			Data_memory[116] <= 32'd0; 
			Data_memory[117] <= 32'd0; 
			Data_memory[118] <= 32'd0; 
			Data_memory[119] <= 32'd0; 
			Data_memory[120] <= 32'd0; 
			Data_memory[121] <= 32'd0; 
			Data_memory[122] <= 32'd0; 
			Data_memory[123] <= 32'd0; 
			Data_memory[124] <= 32'd0; 
			Data_memory[125] <= 32'd0; 
			Data_memory[126] <= 32'd0; 
			Data_memory[127] <= 32'd0;
			$display("RESET MODE");	
		end   	
	
		else
		begin
			Data_memory[0] <=	Data_memory[0]	;
			Data_memory[1] <=	Data_memory[1]	;
			Data_memory[2] <=	Data_memory[2]	;
			Data_memory[3] <=	Data_memory[3]	;
			Data_memory[4] <=	Data_memory[4]	;
			Data_memory[5] <=	Data_memory[5]	;
			Data_memory[6] <=	Data_memory[6]	;
			Data_memory[7] <=	Data_memory[7]	;
			Data_memory[8] <=	Data_memory[8]	;
			Data_memory[9] <=	Data_memory[9]	;
			Data_memory[10] <= 	Data_memory[10]	;
			Data_memory[11] <=	Data_memory[11]	;
			Data_memory[12] <=	Data_memory[12]	;
			Data_memory[13] <=	Data_memory[13]	;
			Data_memory[14] <=	Data_memory[14]	;
			Data_memory[15] <=	Data_memory[15]	;
			Data_memory[16] <=	Data_memory[16]	;
			Data_memory[17] <=	Data_memory[17]	;
			Data_memory[18] <=	Data_memory[18]	;
			Data_memory[19] <=	Data_memory[19]	;
			Data_memory[20] <=	Data_memory[20]	;
			Data_memory[21] <=	Data_memory[21]	;
			Data_memory[22] <=	Data_memory[22]	;
			Data_memory[23] <=	Data_memory[23]	;
			Data_memory[24] <=	Data_memory[24]	;
			Data_memory[25] <=	Data_memory[25]	;
			Data_memory[26] <=	Data_memory[26]	;
			Data_memory[27] <=	Data_memory[27]	;
			Data_memory[28] <=	Data_memory[28]	;
			Data_memory[29] <=	Data_memory[29]	;
			Data_memory[30] <=	Data_memory[30]	;
			Data_memory[31] <=	Data_memory[31]	;
			Data_memory[32] <=	Data_memory[32]	;
			Data_memory[33] <=	Data_memory[33]	;
			Data_memory[34] <=	Data_memory[34]	;
			Data_memory[35] <=	Data_memory[35]	;
			Data_memory[36] <=	Data_memory[36]	;
			Data_memory[37] <=	Data_memory[37]	;
			Data_memory[38] <=	Data_memory[38]	;
			Data_memory[39] <=	Data_memory[39]	;
			Data_memory[40] <=	Data_memory[40]	;
			Data_memory[41] <=	Data_memory[41]	;
			Data_memory[42] <=	Data_memory[42]	;
			Data_memory[43] <=	Data_memory[43]	;
			Data_memory[44] <=	Data_memory[44]	;
			Data_memory[45] <=	Data_memory[45]	;
			Data_memory[46] <=	Data_memory[46]	;
			Data_memory[47] <=	Data_memory[47]	;
			Data_memory[48] <=	Data_memory[48]	;
			Data_memory[49] <=	Data_memory[49]	;
			Data_memory[50] <=	Data_memory[50]	;
			Data_memory[51] <=	Data_memory[51]	;
			Data_memory[52] <=	Data_memory[52]	;
			Data_memory[53] <=	Data_memory[53]	;
			Data_memory[54] <=	Data_memory[54]	;
			Data_memory[55] <=	Data_memory[55]	;
			Data_memory[56] <=	Data_memory[56]	;
			Data_memory[57] <=	Data_memory[57]	;
			Data_memory[58] <=	Data_memory[58]	;
			Data_memory[59] <=	Data_memory[59]	;
			Data_memory[60] <=	Data_memory[60]	;
			Data_memory[61] <=	Data_memory[61]	;
			Data_memory[62] <=	Data_memory[62]	;
			Data_memory[63] <=	Data_memory[63]	;
			Data_memory[64] <=	Data_memory[64]	;
			Data_memory[65] <=	Data_memory[65]	;
			Data_memory[66] <=	Data_memory[66]	;
			Data_memory[67] <=	Data_memory[67]	;
			Data_memory[68] <=	Data_memory[68]	;
			Data_memory[69] <=	Data_memory[69]	;
			Data_memory[70] <=	Data_memory[70]	;
			Data_memory[71] <=	Data_memory[71]	;
			Data_memory[72] <=	Data_memory[72]	;
			Data_memory[73] <=	Data_memory[73]	;
			Data_memory[74] <= 	Data_memory[74]	;
			Data_memory[75] <=	Data_memory[75]	;
			Data_memory[76] <=	Data_memory[76]	;
			Data_memory[77] <=	Data_memory[77]	;
			Data_memory[78] <=	Data_memory[78]	;
			Data_memory[79] <=	Data_memory[79]	;
			Data_memory[80] <=	Data_memory[80]	;
			Data_memory[81] <=	Data_memory[81]	;
			Data_memory[82] <=	Data_memory[82]	;
			Data_memory[83] <=	Data_memory[83]	;
			Data_memory[84] <=	Data_memory[84]	;
			Data_memory[85] <=	Data_memory[85]	;
			Data_memory[86] <=	Data_memory[86]	;
			Data_memory[87] <=	Data_memory[87]	;
			Data_memory[88] <=	Data_memory[88]	;
			Data_memory[89] <=	Data_memory[89]	;
			Data_memory[90] <=	Data_memory[90]	;
			Data_memory[91] <=	Data_memory[91]	;
			Data_memory[92] <=	Data_memory[92]	;
			Data_memory[93] <=	Data_memory[93]	;
			Data_memory[94] <=	Data_memory[94]	;
			Data_memory[95] <=	Data_memory[95]	;
			Data_memory[96] <=	Data_memory[96]	;
			Data_memory[97] <=	Data_memory[97]	;
			Data_memory[98] <=	Data_memory[98]	;
			Data_memory[99] <=	Data_memory[99]	;
			Data_memory[100] <=	Data_memory[100]	;
			Data_memory[101] <=	Data_memory[101]	;
			Data_memory[102] <=	Data_memory[102]	;
			Data_memory[103] <=	Data_memory[103]	;
			Data_memory[104] <=	Data_memory[104]	;
			Data_memory[105] <=	Data_memory[105]	;
			Data_memory[106] <=	Data_memory[106]	;
			Data_memory[107] <=	Data_memory[107]	;
			Data_memory[108] <=	Data_memory[108]	;
			Data_memory[109] <=	Data_memory[109]	;
			Data_memory[110] <=	Data_memory[110]	;
			Data_memory[111] <=	Data_memory[111]	;
			Data_memory[112] <=	Data_memory[112]	;
			Data_memory[113] <=	Data_memory[113]	;
			Data_memory[114] <=	Data_memory[114]	;
			Data_memory[115] <=	Data_memory[115]	;
			Data_memory[116] <=	Data_memory[116]	;
			Data_memory[117] <=	Data_memory[117]	;
			Data_memory[118] <=	Data_memory[118]	;
			Data_memory[119] <=	Data_memory[119]	;
			Data_memory[120] <=	Data_memory[120]	;
			Data_memory[121] <=	Data_memory[121]	;
			Data_memory[122] <=	Data_memory[122]	;
			Data_memory[123] <=	Data_memory[123]	;
			Data_memory[124] <=	Data_memory[124]	;
			Data_memory[125] <=	Data_memory[125]	;
			Data_memory[126] <=	Data_memory[126]	;
			Data_memory[127] <=	Data_memory[127]	;

   			//$display("Data_mem_Address: %d", Address);
			if (MemWrite==1) begin
				Data_memory[Address>>2] <= Write_Data;
				//$display("Write_data: %d", Write_Data);
			end
   			//else if	(MemRead == 1) begin
                		//Read_data <= Data_memory[Address>>2];
				//$display("Read_data: %d", Read_data);
   			//end 
			//else Read_data <= 32'h00000000;
   		end

endmodule
