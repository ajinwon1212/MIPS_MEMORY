module Shift_left_2 (
	input [31:0] Shift_left_2_IN,
	output [31:0] Shift_left_2_OUT
	);

	assign Shift_left_2_OUT = Shift_left_2_IN << 2;

endmodule
